module test(
);

initial begin
    $display("Hello World");
    $finish;
end

endmodule

