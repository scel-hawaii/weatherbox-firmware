module test(
    reset
);

input reset;

initial begin
    $display("Hello World");
    $finish;
end

endmodule

